kcsncohacba
